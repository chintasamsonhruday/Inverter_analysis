
** Generated for: hspiceD
** Generated on: Oct  8 19:27:58 2024
** Design library name: class_project1
** Design cell name: NMOS
** Design view name: schematic


**.TEMP 25.0
**.OPTION
**+    ARTIST=2
**+    INGOLD=2
**+    PARHIER=LOCAL
**+    PSF=2

** Library name: class_project1
** Cell name: NMOS
** View name: schematic
m3 y a vdd vdd pch_svt_mac l=16e-9 nfin=8 w=346e-9 multi=1 nf=1 sa=90e-9 sb=90e-9
.END
