** Generated for: hspiceD
** Generated on: Oct  8 16:34:22 2024
** Design library name: ckt1
** Design cell name: inverter1
** Design view name: schematic


**.TEMP 25.0
**.OPTION
**+    ARTIST=2
**+    INGOLD=2
**+    PARHIER=LOCAL
**+    PSF=2

** Library name: ckt1
** Cell name: inverter1
** View name: schematic
m2 y a gnd gnd nch_svt_mac l=16e-9 nfin=8 w=346e-9 multi=1 nf=1 sa=90e-9 sb=90e-9
m3 y a vdd vdd pch_svt_mac l=16e-9 nfin=8 w=346e-9 multi=1 nf=1 sa=90e-9 sb=90e-9
.END
