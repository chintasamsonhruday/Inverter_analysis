** Generated for: hspiceD
** Generated on: Oct  9 18:43:48 2024
** Design library name: class_project1
** Design cell name: Nmos_inverter
** Design view name: schematic


*.TEMP 25.0
*.OPTION
*+    ARTIST=2
*+    INGOLD=2
*+    PARHIER=LOCAL
*+    PSF=2

** Library name: class_project1
** Cell name: Nmos_inverter
** View name: schematic
m1 vout vin gnd gnd nch_svt_mac l=16e-9 nfin=8 w=346e-9 multi=1 nf=1 sa=90e-9 sb=90e-9
m0 vdd  vdd vout gnd nch_svt_mac l=16e-9 nfin=8 w=346e-9 multi=1 nf=1 sa=90e-9 sb=90e-9
.END
